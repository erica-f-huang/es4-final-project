module top(
        input  clock_in,                
        output HSYNC,                   //go to vga adapter
        output VSYNC,                   //go to vga adapter
        output logic [5:0] rgb,         //go to vga adapter
	output locked                   // leave floating
);


logic intermediate_clk;
logic [9:0] curr_col;
logic [9:0] curr_row;
logic valid;

        mypll u_mypll(
                .clock_in(clock_in),            //in
                .clock_out(intermediate_clk),   //out
                .locked(locked)                 //out
        );

        vga u_vga(
                .clk(intermediate_clk),         //in
                .HSYNC(HSYNC),                  //out
                .VSYNC(VSYNC),                  //out
                .valid(valid),                  //out
                .curr_col(curr_col),            //out
                .curr_row(curr_row)             //out
        );

        screen_gen u_screen_gen(
                .col(curr_col),                 //in
                .row(curr_row),                 //in
                .valid(valid),                  //in
                .rgb(rgb)                       //out
        );





endmodule