// /*MAKES A 0*/

// if ((70 < row) & (row <= 80) |
//     (100 < row) & (row <= 110)) begin
//         rgb = white;
// end else
// if ((80 < row) & (row <= 100)) begin
//         if(((20 < col) & (col <= 30)) | 
//            ((35 < col) & (col <= 45))) begin
//                 rgb = white;
//         end else begin
//                 rgb = black;
//         end
// end else begin
//         rgb = black;    
// end  

// /* MAKES A 0 */ 